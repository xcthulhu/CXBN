use work.common_decs.all;

package write_chanc_decs is
      constant A : natural := write_chan'length; -- number of bits
end package;
