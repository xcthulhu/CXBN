use work.common_decs.all;

package charc_decs is
      constant B : natural := char_size; -- number of bits
end package;
